library ieee;

use ieee.std_logic_1164.all;

entity 32bit_register is
    port(
    );
end 32bit_register;

