library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;


entity datapath is
	port(
		signal clock, clear: in std_logic
	);
end datapath;
